module CalcImmediate(input logic [31:0]instrucao, output logic [63:0]immediate);
logic [63:0]calcImmediate;

calcimm =[11:0]instrucao;

endmodule