`timescale 1ps/1ps

module simulClocks;
logic clk;
logic rst;

meuCpu meuClock(.Clk(clk),.Reset(rst));

   localparam CLKPERIOD = 10000;
   localparam CLKDELAY = CLKPERIOD / 2; 

initial begin
clk=1;
end
always #(CLKDELAY) clk = ~clk;

    initial
    begin
        rst = 1'b0;
        #(CLKPERIOD)
        rst = 1'b1;
        #(CLKPERIOD)
        #(CLKPERIOD)
        rst = 1'b0;       
    end

endmodule